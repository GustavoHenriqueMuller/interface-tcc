library IEEE;
use IEEE.std_logic_1164.all;

entity interface_tcc_backend is
end interface_tcc_backend;

architecture arch_interface_tcc_backend is
end arch_interface_tcc_backend;